module Presets(clk, sel, grid);
	parameter gsr = 20;	//grid size
	parameter gsc = 20;
	parameter addr_len = 8;
	input clk;
	input [2:0] sel;
	output reg [gsr*gsc:0] grid;
	
	wire [addr_len-1:0]hgs_r = 0; //half grid size
	wire [addr_len-1:0]hgs_c = 0;

	wire [gsr*gsc:0] rand;
	Randomizer #(gsr, gsc) (clk, rand);
	
	always @(sel) begin
		grid = 0;
		case (sel)
			0: begin
			end
			1: begin
				//glider
				grid[gsc*(hgs_r+0) + (0+hgs_c)] = 1;
				grid[gsc*(hgs_r+0) + (1+hgs_c)] = 1;
				grid[gsc*(hgs_r+1) + (0+hgs_c)] = 1;
				grid[gsc*(hgs_r+1) + (2+hgs_c)] = 1;
				grid[gsc*(hgs_r+2) + (0+hgs_c)] = 1;
			end
			2: begin
				//pulsar
				grid[gsc*(hgs_r+0) + (3+hgs_c)] = 1;
				grid[gsc*(hgs_r+0) + (4+hgs_c)] = 1; 
				grid[gsc*(hgs_r+0) + (5+hgs_c)] = 1; 
				grid[gsc*(hgs_r+0) + (9+hgs_c)] = 1; 
				grid[gsc*(hgs_r+0) + (10+hgs_c)] = 1;
				grid[gsc*(hgs_r+0) + (11+hgs_c)] = 1;
				grid[gsc*(hgs_r+2) + (1+hgs_c)] = 1; 
				grid[gsc*(hgs_r+2) + (6+hgs_c)] = 1; 
				grid[gsc*(hgs_r+2) + (8+hgs_c)] = 1;
				grid[gsc*(hgs_r+2) + (13+hgs_c)] = 1;
				grid[gsc*(hgs_r+3) + (1+hgs_c)] = 1;
				grid[gsc*(hgs_r+3) + (6+hgs_c)] = 1;
				grid[gsc*(hgs_r+3) + (8+hgs_c)] = 1;
				grid[gsc*(hgs_r+3) + (13+hgs_c)] = 1;
				grid[gsc*(hgs_r+4) + (1+hgs_c)] = 1;
				grid[gsc*(hgs_r+4) + (6+hgs_c)] = 1;
				grid[gsc*(hgs_r+4) + (8+hgs_c)] = 1;
				grid[gsc*(hgs_r+4) + (13+hgs_c)] = 1;
				grid[gsc*(hgs_r+5) + (3+hgs_c)] = 1;
				grid[gsc*(hgs_r+5) + (4+hgs_c)] = 1;
				grid[gsc*(hgs_r+5) + (5+hgs_c)] = 1;
				grid[gsc*(hgs_r+5) + (9+hgs_c)] = 1;
				grid[gsc*(hgs_r+5) + (10+hgs_c)] = 1;
				grid[gsc*(hgs_r+5) + (11+hgs_c)] = 1;
				grid[gsc*(hgs_r+7) + (3+hgs_c)] = 1;
				grid[gsc*(hgs_r+7) + (4+hgs_c)] = 1;
				grid[gsc*(hgs_r+7) + (5+hgs_c)] = 1;
				grid[gsc*(hgs_r+7) + (9+hgs_c)] = 1;
				grid[gsc*(hgs_r+7) + (10+hgs_c)] = 1;
				grid[gsc*(hgs_r+7) + (11+hgs_c)] = 1;
				grid[gsc*(hgs_r+8) + (1+hgs_c)] = 1;
				grid[gsc*(hgs_r+8) + (6+hgs_c)] = 1;
				grid[gsc*(hgs_r+8) + (8+hgs_c)] = 1;
				grid[gsc*(hgs_r+8) + (13+hgs_c)] = 1;
				grid[gsc*(hgs_r+9) + (1+hgs_c)] = 1;
				grid[gsc*(hgs_r+9) + (6+hgs_c)] = 1;
				grid[gsc*(hgs_r+9) + (8+hgs_c)] = 1;
				grid[gsc*(hgs_r+9) + (13+hgs_c)] = 1;
				grid[gsc*(hgs_r+10) + (1+hgs_c)] = 1;
				grid[gsc*(hgs_r+10) + (6+hgs_c)] = 1;
				grid[gsc*(hgs_r+10) + (8+hgs_c)] = 1;
				grid[gsc*(hgs_r+10) + (13+hgs_c)] = 1;
				grid[gsc*(hgs_r+12) + (3+hgs_c)] = 1;
				grid[gsc*(hgs_r+12) + (4+hgs_c)] = 1;
				grid[gsc*(hgs_r+12) + (5+hgs_c)] = 1;
				grid[gsc*(hgs_r+12) + (9+hgs_c)] = 1;
				grid[gsc*(hgs_r+12) + (10+hgs_c)] = 1;
				grid[gsc*(hgs_r+12) + (11+hgs_c)] = 1;
			end
			3: begin
				//lightweight spaceship
				grid[gsc*(hgs_r+0) + (0+hgs_c)] = 1;
				grid[gsc*(hgs_r+0) + (3+hgs_c)] = 1;
				grid[gsc*(hgs_r+1) + (4+hgs_c)] = 1;
				grid[gsc*(hgs_r+2) + (0+hgs_c)] = 1;
				grid[gsc*(hgs_r+2) + (4+hgs_c)] = 1;
				grid[gsc*(hgs_r+3) + (1+hgs_c)] = 1;
				grid[gsc*(hgs_r+3) + (2+hgs_c)] = 1;
				grid[gsc*(hgs_r+3) + (3+hgs_c)] = 1;
				grid[gsc*(hgs_r+3) + (4+hgs_c)] = 1;
			end
			4: begin
				//gosper's glider gun
				grid[gsc*(hgs_r+0) + (24+hgs_c)] = 1;
				grid[gsc*(hgs_r+1) + (22+hgs_c)] = 1;
				grid[gsc*(hgs_r+1) + (24+hgs_c)] = 1;
				grid[gsc*(hgs_r+2) + (12+hgs_c)] = 1;
				grid[gsc*(hgs_r+2) + (13+hgs_c)] = 1;
				grid[gsc*(hgs_r+2) + (20+hgs_c)] = 1;
				grid[gsc*(hgs_r+2) + (21+hgs_c)] = 1;
				grid[gsc*(hgs_r+2) + (34+hgs_c)] = 1;
				grid[gsc*(hgs_r+2) + (35+hgs_c)] = 1;
				grid[gsc*(hgs_r+3) + (11+hgs_c)] = 1;
				grid[gsc*(hgs_r+3) + (15+hgs_c)] = 1;
				grid[gsc*(hgs_r+3) + (20+hgs_c)] = 1;
				grid[gsc*(hgs_r+3) + (21+hgs_c)] = 1;
				grid[gsc*(hgs_r+3) + (34+hgs_c)] = 1;
				grid[gsc*(hgs_r+3) + (35+hgs_c)] = 1;
				grid[gsc*(hgs_r+4) + (0+hgs_c)] = 1;
				grid[gsc*(hgs_r+4) + (1+hgs_c)] = 1;
				grid[gsc*(hgs_r+4) + (10+hgs_c)] = 1;
				grid[gsc*(hgs_r+4) + (16+hgs_c)] = 1;
				grid[gsc*(hgs_r+4) + (20+hgs_c)] = 1;
				grid[gsc*(hgs_r+4) + (21+hgs_c)] = 1;
				grid[gsc*(hgs_r+5) + (0+hgs_c)] = 1;
				grid[gsc*(hgs_r+5) + (1+hgs_c)] = 1;
				grid[gsc*(hgs_r+5) + (10+hgs_c)] = 1;
				grid[gsc*(hgs_r+5) + (14+hgs_c)] = 1;
				grid[gsc*(hgs_r+5) + (16+hgs_c)] = 1;
				grid[gsc*(hgs_r+5) + (17+hgs_c)] = 1;
				grid[gsc*(hgs_r+5) + (22+hgs_c)] = 1;
				grid[gsc*(hgs_r+5) + (24+hgs_c)] = 1;
				grid[gsc*(hgs_r+6) + (10+hgs_c)] = 1;
				grid[gsc*(hgs_r+6) + (16+hgs_c)] = 1;
				grid[gsc*(hgs_r+6) + (24+hgs_c)] = 1;
				grid[gsc*(hgs_r+7) + (11+hgs_c)] = 1;
				grid[gsc*(hgs_r+7) + (15+hgs_c)] = 1;
				grid[gsc*(hgs_r+8) + (12+hgs_c)] = 1;
				grid[gsc*(hgs_r+8) + (13+hgs_c)] = 1;
			end
			5: begin
				grid[gsr*gsc:0] <= rand[gsr*gsc:0];
			end
			default: begin end
		endcase
	end
endmodule

//LFSR-based Randomizer
module Randomizer(clk, grid);
	parameter gsr = 20;	//grid size
	parameter gsc = 20;
	input clk;
	output reg [gsr*gsc:0] grid = 1200'b00110010101110101010111100101101011111110011011100101101111101100000111100000100101110101001110000010111010111010011110100001111100010000000011001100001011111100001011100001001000011110110010000011101010110100001001000010110100011101100010011000110111001100110001100011101001011011101001010001010100001000100010010110111101111101001001100000110111001110001110100010000011010111000111110010110110000111110001100101001111111110111010010111100011110101110010011001111101100101011001000110111001101100010111111111101000011101110000001011110110000100001101100000011101010110000110111010100000010100110001111000101000010100110010110010011101011101010000011101111000101110000000100101111111010000111010011000111100010100101100110110011110000101111011001011110111010010110100001010101111011011001100001011110111110101011110110111000000000111000100100101110001011011011001000110110111011110111011000000000000011001011100100000011000000000011101001101010100101011111010101101010010010110000011100001001100000100011001101010001010001101000000010011011001001010011011111101011001011011001100100100111010100010110000000101000011001000110101100110010000110011111111010010001101100100110100100010010010111001001101000000011000001010000110000100010100100101010101010010010110010111010001110010001011110100010101011001010101010011001011000100101011101011011000001111000001001111111110001001000110000010000000000001111100011101101001101010011010010011000101101000001110000101000001111100100000100111000011101001100011001110110011011110010111011111001110110100100010100010001100101001110110000010110101100011000111011010000000100000001111000101011001101101011001111000100100011010001100010110011111101111101010000110110111010011101000111000110110100001011000010110010101111010111011011110010100110110000001110000000111110001110110101101001111011111001101100000101101110110100011001010011000001000101100101100101000001111010011101110011011110011100000011101000110111011100101010011000000101001000001000001111110011110100001101111111001110110000110000010101011100110010100000100100101110001001011100110111000001001110000110001100111111010101011111001100001110011010010110111000110111100110100000001111111011110101010110001000011101110000011001001111010110000100001111010001100000011011000010010010110101110010000101011110100010101110011111001001000001011010100111110010101010011110011001110000001101010100111110100000000011100001100101101000101100011101101011000011111110010110011100011100111001000011001000101011010010101000111011110101011011011000001000001110001001011101101100101000101101010100100000111010111001010110000011111101110000110110100110010001101001001011011010010110010111000000101101100110001110101101111111101001010101111110100101010101110110011010001111111010000010000111110000100110011111010011100010110011101111100101001011101111111101111000101000111100000111101111101110101001001100000000110100010100000010110001001010010111001011111000011101100100110001011111101001110010110011111010111101110100000101010010001000010001111101001001100111100100010110011011110110111110001101100010111000011111000100111000000111011101001111110001010000001001011010010100101010011100000011000010111011100010101001001010011110000000000110011001010110001011110110000001001010110110001001111010101100110101011000100001100010001011110101000010000011001001011111100101011010111011101010010110000000001101110100000011111011110101010000000100011001000010001110011100100011100100100110110101110001100000101111100011010011111010111010100101101011011001100100101000001011010110011000110111101011101001110101000000011010010010110110001010000001000101101100011100101100001110101000111101001001111000010100001011111100100101111011111110000011100111100100001001110100101010010001011111110001011111111101100000001011000010110111010001011010110110011001101100100010100010101111101001100111110010111110011010110110010101110110111000000110011110010111010010101111011000110101100110100001101000101111100111100111110101000100111011101100011111001100010101011010101000100111010001011101111100010000110100010100110011000101011100100010001000111010010010110010111011011011101000000101011100111011011011001010101001110101110101111110000110000110100111110110011010101000101101000101101111000000010110111100110111011100110111101001100000111000100110100100011110101001101011010010111110010001110111001000010110110101101000011110110110101010010011000111000111011111111101110000101100000110110101100000000101111110110111110001011011011111011011001111011001010010011001110000111110111100111001111110110001000100101110001001011101001010000001001101111011011100110010100101001111110011101000010100110000100000100111111101111011111010001111100010001110110100111001001011001000100010110010100000110111111011011110110101001000001001101101010011010001010000011110000001110110111011111001100000100010111110101111011110010100110111110001100011111010111010101110110110110100011010010100011111101111100111111010100001010101110100001101101011101110000101010100000011011100111001010110111000011011111100110110100001000110110010010111001111000101001110011000111101110111100110010101100100111100001001000101011001000010000100010011010010000100101010000110101111011101100110111101110000101100010001110110100100101111001100101001010011011100100001010100111100100101100101000010001001101111101111110011000111100011100011011110110111010001010111010100101100101101111011101110000101011101100010101100001101010000110110000011101101100100011011010010110101100110100011010011011000100001011000100000100101011001011110111110000101100000111110110101100000000101000010110010010011011111010110110110010100001010010011101100110100000111100011010110011101111110111001000010010111011011010111100010100001101001111010010010111001001000111111110110011100001001000010000100001010101110011001011001110000100101100010110101011110010100011000111000001110000010111011100001001101100111111111111111101010100001001111110011101101000010101000110011100111001011011100000111000010110011011111100110101001000101000110110111111001011110001111100111001000001110101110101111110100000101100101101001010001100000110001011100001001010100000110001101001011100010010110111100101100100001110011110001100001100101110101011100110001110000101000011100100101110001110011111100011101101100000000111001011011100110010010100101101011100011100000001101001000010001010111101011001101001010010100101011011101100100010001011100010100000110011111001011011100100001100001110111001100100101111100011010010111011101001110100110111111110010010001110001110100011010011100001100000000110111011001000010010111000000001010010110111000100101110001010011010100111011110010000011001111011111111000111110110111011100110010111001101100001010111000101000100111001101111011110001101101100111111010011010010011101100000001000000000111110011001111110000001111110111011100011011010110001011010000010100100111011000101000001011111011000011110000101010100000011101111011101110000100111000000000010000100010111000011100100101001111101001100111000100011011101111111011001001011010010100100010111101100000111001101011000101101110001001001111100010101001001100100110001010110011000010000100010010111011111011110111010100001010010011110101111011001010010010100100011110111010111110010000001001000010111110110111111000000110011001101001111111010100101011010100001111011001010001000001111010000010110001101101000001000101110000100100100001010011111010110001010110011001010110011110110000100001100101111111100100101000100010101010001001010011010000011101111100011110101011011111010101000011110000111011100110000100101011010110001000100100011011010001111010101101100000001011001001010101100011111000011000101101111000100101100001011001101011111101110100010001110001100110001111011001000010011111010110110011000010100000011101001111101101111101100011011000111010000011110101010101010010011110001010110000010110110111000111000001111010101010100101011111011010111110111000000110111011010111110100000101011010110011010110010000111001001000001001010000110001100110111111101001100000101110110011110000111101010010111100100111110100111000100010000011110011110001110001110000100100001101011010100000111100110110011101101000111010111000001011001101110011000100100110100001010110000011001110111111000111010010011010001101110101110101000001010100100100101110110110000100010010100010110100110011000011101100000010100100111000011100010010111110000100011011110010010010011001101010110000101101011011011101001001010110110101110110000110000111010011011100110001010110010010110011011001011001011110110110100000100100000001111111110011110101010011101100000011000001111111010110011000100011010001111110001010110110100010000111000111010100000110111100101100000001110111000101101011011111001110000111010010010110110101001101000111011000011111110111001010000010111011101100110110111100100110000000100100011110011101011001011000110110000100101100000010110011000101011100010001111100001100000010100011110110110101011110110100010101110100111101011000111000110100111000001111101001011111101001110111101001001101000111100100011000111011011101111100001011101010111100010111001111111001110010011010010101101010010111110100110010011110100110101101010111110110101001010100110100100011010000101001111110011111001000100011001111111100101010100001111101011000001001101000111011101100110011010101110011101110110011011101010010100101001111111100100011000011100100011100000010011000000011111010000001100000110101100101001110000000111111100000001010110111101011011101110111000110010110010101011111011100111011111110111111010101110110100001110001100011001101101100010010001101010010011101110110001010001000010001111011011111001011010111001100001101011110111100111111010101111001110011111111010011011001001111000101111001000010000110011001110100010100010011010000000101100110111000000110100010110110100000001000011110011000101111010101110010001101000000000101110011000100010000111001101000010111010000100110100110101011110010000010100001111110100101110001100000001110110011101011110100001101110100100010111011001101011000111111101100110110000010101010111101111110100100011111010011010010011111100011001110111111101100011001110110100010011000010000110110010101011011100000111000100000010100100001110111010111000000111010111101001111101000000001111000111000011001001000011110000110010011111111001000100110111110101110000010111101111101110010110010100011101101001011111100011100011100010001001011001111110101101010101011000110100001010111100101110001100000010010111110101001000110000000000100100000111011001100001101011101000101111100101101000100011110111110010011010000101010001110010110100111011100001100000000111011010110001000011101001001001010000001000000111111011111111000001001101001001100110011100110111001100000001010010010110000010011110101100111110001101100000101110011000100001110000111011111111110110111010000001000010010000101101011011010101111101100011111101011011100000001100000010000101110010100101100110001100110110101101100001111011010000111011111001111000010001000001110111001010010000100001011111000000001101111011110101000000100001100001111100101000111000100110110100011001000110011010100111010000110110101010110111001111001010000111100010101000110011111001111100100101110000101011111101000110000111000010111100101110101101001011110100000000000010110010100101100101110000101011100011111110110000010111101011100111000111111001001001100001011110000011001001101110011010110010001100111010110101111100000011000110101110000000100111110100001000011100001011100011111011011101010001111101101101010001101111001001001110001001111101100001111100101111110100111101010111010000111111100101000101011100101111110010001110000010111011001110110001000100010110110010011001100111000100010110110010010001110001100011111010101000010000100001110011001111110000000011001101111000111011010011011011000000000110010001001110110101000111110111101110011001100101101010111011000111011111111110011001010010000001100010010111000101110001000100101011010111001001110001111000111101010;
	
	always @(posedge clk) begin
		grid <= {(grid[0]^grid[2]^grid[4]^grid[6]), grid[gsr*gsc:1]};
	end
endmodule
